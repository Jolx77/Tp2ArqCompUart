module uart_rx #(
    parameter N = 8,  // Number of data bits
    parameter M = 1,  // Number of stop bits
    parameter PARITY_EN = 0,  // Enable parity bit (0: disable, 1: enable)
    parameter BAUD_RATE = 9600,  // Baud rate
    parameter CLK_FREQ = 50000000  // Clock frequency
)(
    input wire clk,
    input wire reset,
    input wire rx,
    output reg [N-1:0] data_out,
    output reg valid
);

    // Calculate the number of clock cycles per bit
    localparam integer CYCLES_PER_BIT = CLK_FREQ / BAUD_RATE;
    localparam integer TICK_COUNTER_WIDTH = $clog2(CYCLES_PER_BIT);
    localparam integer BIT_COUNTER_WIDTH = $clog2(N + M + PARITY_EN);

    // State definitions
    typedef enum reg [2:0] {
        IDLE,
        START,
        DATA,
        PARITY,
        STOP
    } state_t;

    state_t state, next_state;

    // Tick counter
    reg [TICK_COUNTER_WIDTH-1:0] tick_counter;

    // Shift register
    reg [N-1:0] shift_reg;
    reg [BIT_COUNTER_WIDTH-1:0] bit_counter;

    // State machine
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= IDLE;
            tick_counter <= 0;
            bit_counter <= 0;
            shift_reg <= 0;
            valid <= 0;
        end else begin
            state <= next_state;
            if (state == START || state == DATA || state == PARITY || state == STOP) begin
                tick_counter <= tick_counter + 1;
            end else begin
                tick_counter <= 0;
            end
        end
    end

    always @(*) begin
        next_state = state;
        case (state)
            IDLE: begin
                if (rx == 0) begin
                    next_state = START;
                end
            end
            START: begin
                if (tick_counter == (CYCLES_PER_BIT / 2 - 1)) begin
                    next_state = DATA;
                    tick_counter = 0;
                end
            end
            DATA: begin
                if (tick_counter == (CYCLES_PER_BIT - 1)) begin
                    shift_reg = {rx, shift_reg[N-1:1]};
                    bit_counter = bit_counter + 1;
                    tick_counter = 0;
                    if (bit_counter == N-1) begin
                        if (PARITY_EN) begin
                            next_state = PARITY;
                        end else begin
                            next_state = STOP;
                        end
                    end
                end
            end
            PARITY: begin
                if (tick_counter == (CYCLES_PER_BIT - 1)) begin
                    // Handle parity bit if needed
                    next_state = STOP;
                    tick_counter = 0;
                end
            end
            STOP: begin
                if (tick_counter == (CYCLES_PER_BIT - 1)) begin
                    bit_counter = bit_counter + 1;
                    tick_counter = 0;
                    if (bit_counter == M) begin
                        next_state = IDLE;
                        data_out = shift_reg;
                        valid = 1;
                    end
                end
            end
        endcase
    end

endmodule



module uart_tx #(
    parameter N = 8,  // Number of data bits
    parameter M = 1,  // Number of stop bits
    parameter PARITY_EN = 0,  // Enable parity bit (0: disable, 1: enable)
    parameter BAUD_RATE = 9600,  // Baud rate
    parameter CLK_FREQ = 50000000  // Clock frequency
)(
    input wire clk,
    input wire reset,
    input wire start_tx,
    input wire [N-1:0] data_in,
    output reg tx,
    output reg busy
);

    // Calculate the number of clock cycles per bit
    localparam integer CYCLES_PER_BIT = CLK_FREQ / BAUD_RATE;
    localparam integer TICK_COUNTER_WIDTH = $clog2(CYCLES_PER_BIT);
    localparam integer BIT_COUNTER_WIDTH = $clog2(N + M + PARITY_EN);

    // State definitions
    typedef enum reg [2:0] {
        IDLE,
        START,
        DATA,
        PARITY,
        STOP
    } state_t;

    state_t state, next_state;

    // Tick counter
    reg [TICK_COUNTER_WIDTH-1:0] tick_counter;

    // Shift register
    reg [N-1:0] shift_reg;
    reg [BIT_COUNTER_WIDTH-1:0] bit_counter;

    // Parity bit
    reg parity_bit;

    // State machine
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            state <= IDLE;
            tick_counter <= 0;
            bit_counter <= 0;
            shift_reg <= 0;
            parity_bit <= 0;
            tx <= 1;
            busy <= 0;
        end else begin
            state <= next_state;
            if (state == START || state == DATA || state == PARITY || state == STOP) begin
                tick_counter <= tick_counter + 1;
            end else begin
                tick_counter <= 0;
            end
        end
    end

    always @(*) begin
        next_state = state;
        case (state)
            IDLE: begin
                if (start_tx) begin
                    next_state = START;
                    shift_reg = data_in;
                    parity_bit = ^data_in;  // Calculate parity bit
                    busy = 1;
                end
            end
            START: begin
                if (tick_counter == (CYCLES_PER_BIT - 1)) begin
                    next_state = DATA;
                    tick_counter = 0;
                    tx = 0;  // Start bit
                end
            end
            DATA: begin
                if (tick_counter == (CYCLES_PER_BIT - 1)) begin
                    tx = shift_reg[0];
                    shift_reg = shift_reg >> 1;
                    bit_counter = bit_counter + 1;
                    tick_counter = 0;
                    if (bit_counter == N-1) begin
                        if (PARITY_EN) begin
                            next_state = PARITY;
                        end else begin
                            next_state = STOP;
                        end
                    end
                end
            end
            PARITY: begin
                if (tick_counter == (CYCLES_PER_BIT - 1)) begin
                    tx = parity_bit;
                    next_state = STOP;
                    tick_counter = 0;
                end
            end
            STOP: begin
                if (tick_counter == (CYCLES_PER_BIT - 1)) begin
                    tx = 1;  // Stop bit
                    bit_counter = bit_counter + 1;
                    tick_counter = 0;
                    if (bit_counter == M) begin
                        next_state = IDLE;
                        busy = 0;
                    end
                end
            end
        endcase
    end

endmodule

